.TITLE statci_adder
.include components.sp
*Subcircuit of an adder unit
.subckt STAT_FA VDD CI
+P0 P1 P2 P3
+D0 D1 D2 D3
+NG0 NG1 NG2 NG3
+C0 C1 C2 C3
X1 VDD CI P0 D0 NG0 C0 STAT_MC_CHAIN
X2 VDD C0 P1 D1 NG1 C1 STAT_MC_CHAIN
X3 VDD C1 P2 D2 NG2 C2 STAT_MC_CHAIN
X4 VDD C2 P3 D3 NG3 C3 STAT_MC_CHAIN
.ends

*Subcircuit of a 4bit carry bypass adder
.subckt STAT_4BIT VDD A0 A1 A2 A3 B0 B1 B2 B3 CI S0 S1 S2 S3 CO
X1 VDD A0 B0 P0 XOR
X2 VDD A1 B1 P1 XOR
X3 VDD A2 B2 P2 XOR
X4 VDD A3 B3 P3 XOR
X5 VDD A0 B0 NG0 NAND
X6 VDD A1 B1 NG1 NAND
X7 VDD A2 B2 NG2 NAND
X8 VDD A3 B3 NG3 NAND
X9 VDD A0 B0 D0 NOR
X10 VDD A1 B1 D1 NOR
X11 VDD A2 B2 D2 NOR
X12 VDD A3 B3 D3 NOR
X13 VDD CI P0 P1 P2 P3 D0 D1 D2 D3 NG0 NG1 NG2 NG3 C0 C1 C2 C3 STAT_FA
X14 VDD P0 P1 1 NAND
X15 VDD P2 P3 2 NAND
X16 VDD 1 2 SEL NOR
X17 VDD CI C3 SEL CO MUX $If SEL(P0P1P2P3) == 1 bypass CI immediately
X18 VDD P0 CI S0 XOR
X19 VDD P1 C0 S1 XOR
X20 VDD P2 C1 S2 XOR
X21 VDD P3 C2 S3 XOR
.ends

*Subcircuit of a 16bit carry bypass adder
.subckt STAT_16BIT VDD CI CO 
+A0 A1 A2 A3 A4 A5 A6 A7 A8 A9 A10 A11 A12 A13 A14 A15
+B0 B1 B2 B3 B4 B5 B6 B7 B8 B9 B10 B11 B12 B13 B14 B15
+S0 S1 S2 S3 S4 S5 S6 S7 S8 S9 S10 S11 S12 S13 S14 S15
X1 VDD A0 A1 A2 A3 B0 B1 B2 B3 CI S0 S1 S2 S3 CO3 STAT_4BIT
*X11 VDD CO3! NCO3 INV
*X12 VDD NCO3 CO3 INV
X2 VDD A4 A5 A6 A7 B4 B5 B6 B7 CO3 S4 S5 S6 S7 CO7 STAT_4BIT
*X21 VDD CO7! NCO7 INV
*X22 VDD NCO7 CO7 INV
X3 VDD A8 A9 A10 A11 B8 B9 B10 B11 CO7 S8 S9 S10 S11 CO11 STAT_4BIT
*X31 VDD CO11! NCO11 INV
*X32 VDD NCO11 CO11 INV
X4 VDD A12 A13 A14 A15 B12 B13 B14 B15 CO11 S12 S13 S14 S15 CO STAT_4BIT
*X41 VDD CO! NCO INV
*X42 VDD NCO CO INV
.ends

*****CRITICAL PATH DELAY*****
V1 vd 0 DC=3.3
V2 vclk 0 PULSE(0 3.3 50ns 1ns 1ns 100ns 202ns)


X1 vd 0 cout
+vd vd vd vd vd vd vd vd vd vd vd vd vd vd vd 0 
+vclk 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0
+S0 S1 S2 S3 S4 S5 S6 S7 S8 S9 S10 S11 S12 S13 S14 S15 STAT_16BIT

.tran 1ns 1000ns 
.MEASURE TRAN tdlay_CO TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(cout) VAL=1.65 RISE = 1

.MEASURE TRAN tdlay_S0 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S0) VAL=1.65 CROSS = 1

.MEASURE TRAN tdlay_S1 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S1) VAL=1.65 CROSS = 1

.MEASURE TRAN tdlay_S2 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S2) VAL=1.65 CROSS = 1

.MEASURE TRAN tdlay_S3 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S3) VAL=1.65 CROSS = 1

.MEASURE TRAN tdlay_S4 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S4) VAL=1.65 CROSS = 1

.MEASURE TRAN tdlay_S5 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S5) VAL=1.65 CROSS = 1

.MEASURE TRAN tdlay_S6 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S6) VAL=1.65 CROSS = 1

.MEASURE TRAN tdlay_S7 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S7) VAL=1.65 CROSS = 1

.MEASURE TRAN tdlay_S8 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S8) VAL=1.65 CROSS = 1

.MEASURE TRAN tdlay_S9 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S9) VAL=1.65 CROSS = 1

.MEASURE TRAN tdlay_S10 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S10) VAL=1.65 CROSS = 1

.MEASURE TRAN tdlay_S11 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S11) VAL=1.65 CROSS = 1

.MEASURE TRAN tdlay_S12 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S12) VAL=1.65 CROSS = 1

.MEASURE TRAN tdlay_S13 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S13) VAL=1.65 CROSS = 1

.MEASURE TRAN tdlay_S14 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S14) VAL=1.65 CROSS = 1

.MEASURE TRAN tdlay_S15 TRIG V(vclk) VAL = 1.65 RISE=1  
+ TARG V(S15) VAL=1.65 CROSS = 1



.END
